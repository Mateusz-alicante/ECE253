//part 2
module part2(A, B, Function, ALUout);
endmodule
