//part 2
